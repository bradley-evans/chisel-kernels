module VecMul( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [15:0] io_A_0, // @[:@6.4]
  input  [15:0] io_A_1, // @[:@6.4]
  input  [15:0] io_A_2, // @[:@6.4]
  input  [15:0] io_A_3, // @[:@6.4]
  input  [15:0] io_A_4, // @[:@6.4]
  input  [15:0] io_A_5, // @[:@6.4]
  input  [15:0] io_A_6, // @[:@6.4]
  input  [15:0] io_A_7, // @[:@6.4]
  input  [15:0] io_A_8, // @[:@6.4]
  input  [15:0] io_A_9, // @[:@6.4]
  input  [15:0] io_A_10, // @[:@6.4]
  input  [15:0] io_A_11, // @[:@6.4]
  input  [15:0] io_A_12, // @[:@6.4]
  input  [15:0] io_A_13, // @[:@6.4]
  input  [15:0] io_A_14, // @[:@6.4]
  input  [15:0] io_A_15, // @[:@6.4]
  input  [15:0] io_B_0, // @[:@6.4]
  input  [15:0] io_B_1, // @[:@6.4]
  input  [15:0] io_B_2, // @[:@6.4]
  input  [15:0] io_B_3, // @[:@6.4]
  input  [15:0] io_B_4, // @[:@6.4]
  input  [15:0] io_B_5, // @[:@6.4]
  input  [15:0] io_B_6, // @[:@6.4]
  input  [15:0] io_B_7, // @[:@6.4]
  input  [15:0] io_B_8, // @[:@6.4]
  input  [15:0] io_B_9, // @[:@6.4]
  input  [15:0] io_B_10, // @[:@6.4]
  input  [15:0] io_B_11, // @[:@6.4]
  input  [15:0] io_B_12, // @[:@6.4]
  input  [15:0] io_B_13, // @[:@6.4]
  input  [15:0] io_B_14, // @[:@6.4]
  input  [15:0] io_B_15, // @[:@6.4]
  output [15:0] io_C_0, // @[:@6.4]
  output [15:0] io_C_1, // @[:@6.4]
  output [15:0] io_C_2, // @[:@6.4]
  output [15:0] io_C_3, // @[:@6.4]
  output [15:0] io_C_4, // @[:@6.4]
  output [15:0] io_C_5, // @[:@6.4]
  output [15:0] io_C_6, // @[:@6.4]
  output [15:0] io_C_7, // @[:@6.4]
  output [15:0] io_C_8, // @[:@6.4]
  output [15:0] io_C_9, // @[:@6.4]
  output [15:0] io_C_10, // @[:@6.4]
  output [15:0] io_C_11, // @[:@6.4]
  output [15:0] io_C_12, // @[:@6.4]
  output [15:0] io_C_13, // @[:@6.4]
  output [15:0] io_C_14, // @[:@6.4]
  output [15:0] io_C_15, // @[:@6.4]
  input         io_load, // @[:@6.4]
  output        io_valid // @[:@6.4]
);
  wire [31:0] _T_153; // @[VecMul.scala 42:35:@9.6]
  wire [32:0] _T_154; // @[VecMul.scala 42:21:@10.6]
  wire [31:0] _T_155; // @[VecMul.scala 42:21:@11.6]
  wire [31:0] _T_156; // @[VecMul.scala 42:35:@12.6]
  wire [32:0] _T_157; // @[VecMul.scala 42:21:@13.6]
  wire [31:0] _T_158; // @[VecMul.scala 42:21:@14.6]
  wire [31:0] _T_159; // @[VecMul.scala 42:35:@15.6]
  wire [32:0] _T_160; // @[VecMul.scala 42:21:@16.6]
  wire [31:0] _T_161; // @[VecMul.scala 42:21:@17.6]
  wire [31:0] _T_162; // @[VecMul.scala 42:35:@18.6]
  wire [32:0] _T_163; // @[VecMul.scala 42:21:@19.6]
  wire [31:0] ans_0; // @[VecMul.scala 42:21:@20.6]
  wire [31:0] _T_165; // @[VecMul.scala 42:35:@21.6]
  wire [32:0] _T_166; // @[VecMul.scala 42:21:@22.6]
  wire [31:0] _T_167; // @[VecMul.scala 42:21:@23.6]
  wire [31:0] _T_168; // @[VecMul.scala 42:35:@24.6]
  wire [32:0] _T_169; // @[VecMul.scala 42:21:@25.6]
  wire [31:0] _T_170; // @[VecMul.scala 42:21:@26.6]
  wire [31:0] _T_171; // @[VecMul.scala 42:35:@27.6]
  wire [32:0] _T_172; // @[VecMul.scala 42:21:@28.6]
  wire [31:0] _T_173; // @[VecMul.scala 42:21:@29.6]
  wire [31:0] _T_174; // @[VecMul.scala 42:35:@30.6]
  wire [32:0] _T_175; // @[VecMul.scala 42:21:@31.6]
  wire [31:0] ans_1; // @[VecMul.scala 42:21:@32.6]
  wire [31:0] _T_177; // @[VecMul.scala 42:35:@33.6]
  wire [32:0] _T_178; // @[VecMul.scala 42:21:@34.6]
  wire [31:0] _T_179; // @[VecMul.scala 42:21:@35.6]
  wire [31:0] _T_180; // @[VecMul.scala 42:35:@36.6]
  wire [32:0] _T_181; // @[VecMul.scala 42:21:@37.6]
  wire [31:0] _T_182; // @[VecMul.scala 42:21:@38.6]
  wire [31:0] _T_183; // @[VecMul.scala 42:35:@39.6]
  wire [32:0] _T_184; // @[VecMul.scala 42:21:@40.6]
  wire [31:0] _T_185; // @[VecMul.scala 42:21:@41.6]
  wire [31:0] _T_186; // @[VecMul.scala 42:35:@42.6]
  wire [32:0] _T_187; // @[VecMul.scala 42:21:@43.6]
  wire [31:0] ans_2; // @[VecMul.scala 42:21:@44.6]
  wire [31:0] _T_189; // @[VecMul.scala 42:35:@45.6]
  wire [32:0] _T_190; // @[VecMul.scala 42:21:@46.6]
  wire [31:0] _T_191; // @[VecMul.scala 42:21:@47.6]
  wire [31:0] _T_192; // @[VecMul.scala 42:35:@48.6]
  wire [32:0] _T_193; // @[VecMul.scala 42:21:@49.6]
  wire [31:0] _T_194; // @[VecMul.scala 42:21:@50.6]
  wire [31:0] _T_195; // @[VecMul.scala 42:35:@51.6]
  wire [32:0] _T_196; // @[VecMul.scala 42:21:@52.6]
  wire [31:0] _T_197; // @[VecMul.scala 42:21:@53.6]
  wire [31:0] _T_198; // @[VecMul.scala 42:35:@54.6]
  wire [32:0] _T_199; // @[VecMul.scala 42:21:@55.6]
  wire [31:0] ans_3; // @[VecMul.scala 42:21:@56.6]
  wire [31:0] _T_201; // @[VecMul.scala 42:35:@57.6]
  wire [32:0] _T_202; // @[VecMul.scala 42:21:@58.6]
  wire [31:0] _T_203; // @[VecMul.scala 42:21:@59.6]
  wire [31:0] _T_204; // @[VecMul.scala 42:35:@60.6]
  wire [32:0] _T_205; // @[VecMul.scala 42:21:@61.6]
  wire [31:0] _T_206; // @[VecMul.scala 42:21:@62.6]
  wire [31:0] _T_207; // @[VecMul.scala 42:35:@63.6]
  wire [32:0] _T_208; // @[VecMul.scala 42:21:@64.6]
  wire [31:0] _T_209; // @[VecMul.scala 42:21:@65.6]
  wire [31:0] _T_210; // @[VecMul.scala 42:35:@66.6]
  wire [32:0] _T_211; // @[VecMul.scala 42:21:@67.6]
  wire [31:0] ans_4; // @[VecMul.scala 42:21:@68.6]
  wire [31:0] _T_213; // @[VecMul.scala 42:35:@69.6]
  wire [32:0] _T_214; // @[VecMul.scala 42:21:@70.6]
  wire [31:0] _T_215; // @[VecMul.scala 42:21:@71.6]
  wire [31:0] _T_216; // @[VecMul.scala 42:35:@72.6]
  wire [32:0] _T_217; // @[VecMul.scala 42:21:@73.6]
  wire [31:0] _T_218; // @[VecMul.scala 42:21:@74.6]
  wire [31:0] _T_219; // @[VecMul.scala 42:35:@75.6]
  wire [32:0] _T_220; // @[VecMul.scala 42:21:@76.6]
  wire [31:0] _T_221; // @[VecMul.scala 42:21:@77.6]
  wire [31:0] _T_222; // @[VecMul.scala 42:35:@78.6]
  wire [32:0] _T_223; // @[VecMul.scala 42:21:@79.6]
  wire [31:0] ans_5; // @[VecMul.scala 42:21:@80.6]
  wire [31:0] _T_225; // @[VecMul.scala 42:35:@81.6]
  wire [32:0] _T_226; // @[VecMul.scala 42:21:@82.6]
  wire [31:0] _T_227; // @[VecMul.scala 42:21:@83.6]
  wire [31:0] _T_228; // @[VecMul.scala 42:35:@84.6]
  wire [32:0] _T_229; // @[VecMul.scala 42:21:@85.6]
  wire [31:0] _T_230; // @[VecMul.scala 42:21:@86.6]
  wire [31:0] _T_231; // @[VecMul.scala 42:35:@87.6]
  wire [32:0] _T_232; // @[VecMul.scala 42:21:@88.6]
  wire [31:0] _T_233; // @[VecMul.scala 42:21:@89.6]
  wire [31:0] _T_234; // @[VecMul.scala 42:35:@90.6]
  wire [32:0] _T_235; // @[VecMul.scala 42:21:@91.6]
  wire [31:0] ans_6; // @[VecMul.scala 42:21:@92.6]
  wire [31:0] _T_237; // @[VecMul.scala 42:35:@93.6]
  wire [32:0] _T_238; // @[VecMul.scala 42:21:@94.6]
  wire [31:0] _T_239; // @[VecMul.scala 42:21:@95.6]
  wire [31:0] _T_240; // @[VecMul.scala 42:35:@96.6]
  wire [32:0] _T_241; // @[VecMul.scala 42:21:@97.6]
  wire [31:0] _T_242; // @[VecMul.scala 42:21:@98.6]
  wire [31:0] _T_243; // @[VecMul.scala 42:35:@99.6]
  wire [32:0] _T_244; // @[VecMul.scala 42:21:@100.6]
  wire [31:0] _T_245; // @[VecMul.scala 42:21:@101.6]
  wire [31:0] _T_246; // @[VecMul.scala 42:35:@102.6]
  wire [32:0] _T_247; // @[VecMul.scala 42:21:@103.6]
  wire [31:0] ans_7; // @[VecMul.scala 42:21:@104.6]
  wire [31:0] _T_249; // @[VecMul.scala 42:35:@105.6]
  wire [32:0] _T_250; // @[VecMul.scala 42:21:@106.6]
  wire [31:0] _T_251; // @[VecMul.scala 42:21:@107.6]
  wire [31:0] _T_252; // @[VecMul.scala 42:35:@108.6]
  wire [32:0] _T_253; // @[VecMul.scala 42:21:@109.6]
  wire [31:0] _T_254; // @[VecMul.scala 42:21:@110.6]
  wire [31:0] _T_255; // @[VecMul.scala 42:35:@111.6]
  wire [32:0] _T_256; // @[VecMul.scala 42:21:@112.6]
  wire [31:0] _T_257; // @[VecMul.scala 42:21:@113.6]
  wire [31:0] _T_258; // @[VecMul.scala 42:35:@114.6]
  wire [32:0] _T_259; // @[VecMul.scala 42:21:@115.6]
  wire [31:0] ans_8; // @[VecMul.scala 42:21:@116.6]
  wire [31:0] _T_261; // @[VecMul.scala 42:35:@117.6]
  wire [32:0] _T_262; // @[VecMul.scala 42:21:@118.6]
  wire [31:0] _T_263; // @[VecMul.scala 42:21:@119.6]
  wire [31:0] _T_264; // @[VecMul.scala 42:35:@120.6]
  wire [32:0] _T_265; // @[VecMul.scala 42:21:@121.6]
  wire [31:0] _T_266; // @[VecMul.scala 42:21:@122.6]
  wire [31:0] _T_267; // @[VecMul.scala 42:35:@123.6]
  wire [32:0] _T_268; // @[VecMul.scala 42:21:@124.6]
  wire [31:0] _T_269; // @[VecMul.scala 42:21:@125.6]
  wire [31:0] _T_270; // @[VecMul.scala 42:35:@126.6]
  wire [32:0] _T_271; // @[VecMul.scala 42:21:@127.6]
  wire [31:0] ans_9; // @[VecMul.scala 42:21:@128.6]
  wire [31:0] _T_273; // @[VecMul.scala 42:35:@129.6]
  wire [32:0] _T_274; // @[VecMul.scala 42:21:@130.6]
  wire [31:0] _T_275; // @[VecMul.scala 42:21:@131.6]
  wire [31:0] _T_276; // @[VecMul.scala 42:35:@132.6]
  wire [32:0] _T_277; // @[VecMul.scala 42:21:@133.6]
  wire [31:0] _T_278; // @[VecMul.scala 42:21:@134.6]
  wire [31:0] _T_279; // @[VecMul.scala 42:35:@135.6]
  wire [32:0] _T_280; // @[VecMul.scala 42:21:@136.6]
  wire [31:0] _T_281; // @[VecMul.scala 42:21:@137.6]
  wire [31:0] _T_282; // @[VecMul.scala 42:35:@138.6]
  wire [32:0] _T_283; // @[VecMul.scala 42:21:@139.6]
  wire [31:0] ans_10; // @[VecMul.scala 42:21:@140.6]
  wire [31:0] _T_285; // @[VecMul.scala 42:35:@141.6]
  wire [32:0] _T_286; // @[VecMul.scala 42:21:@142.6]
  wire [31:0] _T_287; // @[VecMul.scala 42:21:@143.6]
  wire [31:0] _T_288; // @[VecMul.scala 42:35:@144.6]
  wire [32:0] _T_289; // @[VecMul.scala 42:21:@145.6]
  wire [31:0] _T_290; // @[VecMul.scala 42:21:@146.6]
  wire [31:0] _T_291; // @[VecMul.scala 42:35:@147.6]
  wire [32:0] _T_292; // @[VecMul.scala 42:21:@148.6]
  wire [31:0] _T_293; // @[VecMul.scala 42:21:@149.6]
  wire [31:0] _T_294; // @[VecMul.scala 42:35:@150.6]
  wire [32:0] _T_295; // @[VecMul.scala 42:21:@151.6]
  wire [31:0] ans_11; // @[VecMul.scala 42:21:@152.6]
  wire [31:0] _T_297; // @[VecMul.scala 42:35:@153.6]
  wire [32:0] _T_298; // @[VecMul.scala 42:21:@154.6]
  wire [31:0] _T_299; // @[VecMul.scala 42:21:@155.6]
  wire [31:0] _T_300; // @[VecMul.scala 42:35:@156.6]
  wire [32:0] _T_301; // @[VecMul.scala 42:21:@157.6]
  wire [31:0] _T_302; // @[VecMul.scala 42:21:@158.6]
  wire [31:0] _T_303; // @[VecMul.scala 42:35:@159.6]
  wire [32:0] _T_304; // @[VecMul.scala 42:21:@160.6]
  wire [31:0] _T_305; // @[VecMul.scala 42:21:@161.6]
  wire [31:0] _T_306; // @[VecMul.scala 42:35:@162.6]
  wire [32:0] _T_307; // @[VecMul.scala 42:21:@163.6]
  wire [31:0] ans_12; // @[VecMul.scala 42:21:@164.6]
  wire [31:0] _T_309; // @[VecMul.scala 42:35:@165.6]
  wire [32:0] _T_310; // @[VecMul.scala 42:21:@166.6]
  wire [31:0] _T_311; // @[VecMul.scala 42:21:@167.6]
  wire [31:0] _T_312; // @[VecMul.scala 42:35:@168.6]
  wire [32:0] _T_313; // @[VecMul.scala 42:21:@169.6]
  wire [31:0] _T_314; // @[VecMul.scala 42:21:@170.6]
  wire [31:0] _T_315; // @[VecMul.scala 42:35:@171.6]
  wire [32:0] _T_316; // @[VecMul.scala 42:21:@172.6]
  wire [31:0] _T_317; // @[VecMul.scala 42:21:@173.6]
  wire [31:0] _T_318; // @[VecMul.scala 42:35:@174.6]
  wire [32:0] _T_319; // @[VecMul.scala 42:21:@175.6]
  wire [31:0] ans_13; // @[VecMul.scala 42:21:@176.6]
  wire [31:0] _T_321; // @[VecMul.scala 42:35:@177.6]
  wire [32:0] _T_322; // @[VecMul.scala 42:21:@178.6]
  wire [31:0] _T_323; // @[VecMul.scala 42:21:@179.6]
  wire [31:0] _T_324; // @[VecMul.scala 42:35:@180.6]
  wire [32:0] _T_325; // @[VecMul.scala 42:21:@181.6]
  wire [31:0] _T_326; // @[VecMul.scala 42:21:@182.6]
  wire [31:0] _T_327; // @[VecMul.scala 42:35:@183.6]
  wire [32:0] _T_328; // @[VecMul.scala 42:21:@184.6]
  wire [31:0] _T_329; // @[VecMul.scala 42:21:@185.6]
  wire [31:0] _T_330; // @[VecMul.scala 42:35:@186.6]
  wire [32:0] _T_331; // @[VecMul.scala 42:21:@187.6]
  wire [31:0] ans_14; // @[VecMul.scala 42:21:@188.6]
  wire [31:0] _T_333; // @[VecMul.scala 42:35:@189.6]
  wire [32:0] _T_334; // @[VecMul.scala 42:21:@190.6]
  wire [31:0] _T_335; // @[VecMul.scala 42:21:@191.6]
  wire [31:0] _T_336; // @[VecMul.scala 42:35:@192.6]
  wire [32:0] _T_337; // @[VecMul.scala 42:21:@193.6]
  wire [31:0] _T_338; // @[VecMul.scala 42:21:@194.6]
  wire [31:0] _T_339; // @[VecMul.scala 42:35:@195.6]
  wire [32:0] _T_340; // @[VecMul.scala 42:21:@196.6]
  wire [31:0] _T_341; // @[VecMul.scala 42:21:@197.6]
  wire [31:0] _T_342; // @[VecMul.scala 42:35:@198.6]
  wire [32:0] _T_343; // @[VecMul.scala 42:21:@199.6]
  wire [31:0] ans_15; // @[VecMul.scala 42:21:@200.6]
  assign _T_153 = io_A_0 * io_B_0; // @[VecMul.scala 42:35:@9.6]
  assign _T_154 = {{1'd0}, _T_153}; // @[VecMul.scala 42:21:@10.6]
  assign _T_155 = _T_154[31:0]; // @[VecMul.scala 42:21:@11.6]
  assign _T_156 = io_A_1 * io_B_4; // @[VecMul.scala 42:35:@12.6]
  assign _T_157 = _T_155 + _T_156; // @[VecMul.scala 42:21:@13.6]
  assign _T_158 = _T_155 + _T_156; // @[VecMul.scala 42:21:@14.6]
  assign _T_159 = io_A_2 * io_B_8; // @[VecMul.scala 42:35:@15.6]
  assign _T_160 = _T_158 + _T_159; // @[VecMul.scala 42:21:@16.6]
  assign _T_161 = _T_158 + _T_159; // @[VecMul.scala 42:21:@17.6]
  assign _T_162 = io_A_3 * io_B_12; // @[VecMul.scala 42:35:@18.6]
  assign _T_163 = _T_161 + _T_162; // @[VecMul.scala 42:21:@19.6]
  assign ans_0 = _T_161 + _T_162; // @[VecMul.scala 42:21:@20.6]
  assign _T_165 = io_A_0 * io_B_1; // @[VecMul.scala 42:35:@21.6]
  assign _T_166 = {{1'd0}, _T_165}; // @[VecMul.scala 42:21:@22.6]
  assign _T_167 = _T_166[31:0]; // @[VecMul.scala 42:21:@23.6]
  assign _T_168 = io_A_1 * io_B_5; // @[VecMul.scala 42:35:@24.6]
  assign _T_169 = _T_167 + _T_168; // @[VecMul.scala 42:21:@25.6]
  assign _T_170 = _T_167 + _T_168; // @[VecMul.scala 42:21:@26.6]
  assign _T_171 = io_A_2 * io_B_9; // @[VecMul.scala 42:35:@27.6]
  assign _T_172 = _T_170 + _T_171; // @[VecMul.scala 42:21:@28.6]
  assign _T_173 = _T_170 + _T_171; // @[VecMul.scala 42:21:@29.6]
  assign _T_174 = io_A_3 * io_B_13; // @[VecMul.scala 42:35:@30.6]
  assign _T_175 = _T_173 + _T_174; // @[VecMul.scala 42:21:@31.6]
  assign ans_1 = _T_173 + _T_174; // @[VecMul.scala 42:21:@32.6]
  assign _T_177 = io_A_0 * io_B_2; // @[VecMul.scala 42:35:@33.6]
  assign _T_178 = {{1'd0}, _T_177}; // @[VecMul.scala 42:21:@34.6]
  assign _T_179 = _T_178[31:0]; // @[VecMul.scala 42:21:@35.6]
  assign _T_180 = io_A_1 * io_B_6; // @[VecMul.scala 42:35:@36.6]
  assign _T_181 = _T_179 + _T_180; // @[VecMul.scala 42:21:@37.6]
  assign _T_182 = _T_179 + _T_180; // @[VecMul.scala 42:21:@38.6]
  assign _T_183 = io_A_2 * io_B_10; // @[VecMul.scala 42:35:@39.6]
  assign _T_184 = _T_182 + _T_183; // @[VecMul.scala 42:21:@40.6]
  assign _T_185 = _T_182 + _T_183; // @[VecMul.scala 42:21:@41.6]
  assign _T_186 = io_A_3 * io_B_14; // @[VecMul.scala 42:35:@42.6]
  assign _T_187 = _T_185 + _T_186; // @[VecMul.scala 42:21:@43.6]
  assign ans_2 = _T_185 + _T_186; // @[VecMul.scala 42:21:@44.6]
  assign _T_189 = io_A_0 * io_B_3; // @[VecMul.scala 42:35:@45.6]
  assign _T_190 = {{1'd0}, _T_189}; // @[VecMul.scala 42:21:@46.6]
  assign _T_191 = _T_190[31:0]; // @[VecMul.scala 42:21:@47.6]
  assign _T_192 = io_A_1 * io_B_7; // @[VecMul.scala 42:35:@48.6]
  assign _T_193 = _T_191 + _T_192; // @[VecMul.scala 42:21:@49.6]
  assign _T_194 = _T_191 + _T_192; // @[VecMul.scala 42:21:@50.6]
  assign _T_195 = io_A_2 * io_B_11; // @[VecMul.scala 42:35:@51.6]
  assign _T_196 = _T_194 + _T_195; // @[VecMul.scala 42:21:@52.6]
  assign _T_197 = _T_194 + _T_195; // @[VecMul.scala 42:21:@53.6]
  assign _T_198 = io_A_3 * io_B_15; // @[VecMul.scala 42:35:@54.6]
  assign _T_199 = _T_197 + _T_198; // @[VecMul.scala 42:21:@55.6]
  assign ans_3 = _T_197 + _T_198; // @[VecMul.scala 42:21:@56.6]
  assign _T_201 = io_A_4 * io_B_0; // @[VecMul.scala 42:35:@57.6]
  assign _T_202 = {{1'd0}, _T_201}; // @[VecMul.scala 42:21:@58.6]
  assign _T_203 = _T_202[31:0]; // @[VecMul.scala 42:21:@59.6]
  assign _T_204 = io_A_5 * io_B_4; // @[VecMul.scala 42:35:@60.6]
  assign _T_205 = _T_203 + _T_204; // @[VecMul.scala 42:21:@61.6]
  assign _T_206 = _T_203 + _T_204; // @[VecMul.scala 42:21:@62.6]
  assign _T_207 = io_A_6 * io_B_8; // @[VecMul.scala 42:35:@63.6]
  assign _T_208 = _T_206 + _T_207; // @[VecMul.scala 42:21:@64.6]
  assign _T_209 = _T_206 + _T_207; // @[VecMul.scala 42:21:@65.6]
  assign _T_210 = io_A_7 * io_B_12; // @[VecMul.scala 42:35:@66.6]
  assign _T_211 = _T_209 + _T_210; // @[VecMul.scala 42:21:@67.6]
  assign ans_4 = _T_209 + _T_210; // @[VecMul.scala 42:21:@68.6]
  assign _T_213 = io_A_4 * io_B_1; // @[VecMul.scala 42:35:@69.6]
  assign _T_214 = {{1'd0}, _T_213}; // @[VecMul.scala 42:21:@70.6]
  assign _T_215 = _T_214[31:0]; // @[VecMul.scala 42:21:@71.6]
  assign _T_216 = io_A_5 * io_B_5; // @[VecMul.scala 42:35:@72.6]
  assign _T_217 = _T_215 + _T_216; // @[VecMul.scala 42:21:@73.6]
  assign _T_218 = _T_215 + _T_216; // @[VecMul.scala 42:21:@74.6]
  assign _T_219 = io_A_6 * io_B_9; // @[VecMul.scala 42:35:@75.6]
  assign _T_220 = _T_218 + _T_219; // @[VecMul.scala 42:21:@76.6]
  assign _T_221 = _T_218 + _T_219; // @[VecMul.scala 42:21:@77.6]
  assign _T_222 = io_A_7 * io_B_13; // @[VecMul.scala 42:35:@78.6]
  assign _T_223 = _T_221 + _T_222; // @[VecMul.scala 42:21:@79.6]
  assign ans_5 = _T_221 + _T_222; // @[VecMul.scala 42:21:@80.6]
  assign _T_225 = io_A_4 * io_B_2; // @[VecMul.scala 42:35:@81.6]
  assign _T_226 = {{1'd0}, _T_225}; // @[VecMul.scala 42:21:@82.6]
  assign _T_227 = _T_226[31:0]; // @[VecMul.scala 42:21:@83.6]
  assign _T_228 = io_A_5 * io_B_6; // @[VecMul.scala 42:35:@84.6]
  assign _T_229 = _T_227 + _T_228; // @[VecMul.scala 42:21:@85.6]
  assign _T_230 = _T_227 + _T_228; // @[VecMul.scala 42:21:@86.6]
  assign _T_231 = io_A_6 * io_B_10; // @[VecMul.scala 42:35:@87.6]
  assign _T_232 = _T_230 + _T_231; // @[VecMul.scala 42:21:@88.6]
  assign _T_233 = _T_230 + _T_231; // @[VecMul.scala 42:21:@89.6]
  assign _T_234 = io_A_7 * io_B_14; // @[VecMul.scala 42:35:@90.6]
  assign _T_235 = _T_233 + _T_234; // @[VecMul.scala 42:21:@91.6]
  assign ans_6 = _T_233 + _T_234; // @[VecMul.scala 42:21:@92.6]
  assign _T_237 = io_A_4 * io_B_3; // @[VecMul.scala 42:35:@93.6]
  assign _T_238 = {{1'd0}, _T_237}; // @[VecMul.scala 42:21:@94.6]
  assign _T_239 = _T_238[31:0]; // @[VecMul.scala 42:21:@95.6]
  assign _T_240 = io_A_5 * io_B_7; // @[VecMul.scala 42:35:@96.6]
  assign _T_241 = _T_239 + _T_240; // @[VecMul.scala 42:21:@97.6]
  assign _T_242 = _T_239 + _T_240; // @[VecMul.scala 42:21:@98.6]
  assign _T_243 = io_A_6 * io_B_11; // @[VecMul.scala 42:35:@99.6]
  assign _T_244 = _T_242 + _T_243; // @[VecMul.scala 42:21:@100.6]
  assign _T_245 = _T_242 + _T_243; // @[VecMul.scala 42:21:@101.6]
  assign _T_246 = io_A_7 * io_B_15; // @[VecMul.scala 42:35:@102.6]
  assign _T_247 = _T_245 + _T_246; // @[VecMul.scala 42:21:@103.6]
  assign ans_7 = _T_245 + _T_246; // @[VecMul.scala 42:21:@104.6]
  assign _T_249 = io_A_8 * io_B_0; // @[VecMul.scala 42:35:@105.6]
  assign _T_250 = {{1'd0}, _T_249}; // @[VecMul.scala 42:21:@106.6]
  assign _T_251 = _T_250[31:0]; // @[VecMul.scala 42:21:@107.6]
  assign _T_252 = io_A_9 * io_B_4; // @[VecMul.scala 42:35:@108.6]
  assign _T_253 = _T_251 + _T_252; // @[VecMul.scala 42:21:@109.6]
  assign _T_254 = _T_251 + _T_252; // @[VecMul.scala 42:21:@110.6]
  assign _T_255 = io_A_10 * io_B_8; // @[VecMul.scala 42:35:@111.6]
  assign _T_256 = _T_254 + _T_255; // @[VecMul.scala 42:21:@112.6]
  assign _T_257 = _T_254 + _T_255; // @[VecMul.scala 42:21:@113.6]
  assign _T_258 = io_A_11 * io_B_12; // @[VecMul.scala 42:35:@114.6]
  assign _T_259 = _T_257 + _T_258; // @[VecMul.scala 42:21:@115.6]
  assign ans_8 = _T_257 + _T_258; // @[VecMul.scala 42:21:@116.6]
  assign _T_261 = io_A_8 * io_B_1; // @[VecMul.scala 42:35:@117.6]
  assign _T_262 = {{1'd0}, _T_261}; // @[VecMul.scala 42:21:@118.6]
  assign _T_263 = _T_262[31:0]; // @[VecMul.scala 42:21:@119.6]
  assign _T_264 = io_A_9 * io_B_5; // @[VecMul.scala 42:35:@120.6]
  assign _T_265 = _T_263 + _T_264; // @[VecMul.scala 42:21:@121.6]
  assign _T_266 = _T_263 + _T_264; // @[VecMul.scala 42:21:@122.6]
  assign _T_267 = io_A_10 * io_B_9; // @[VecMul.scala 42:35:@123.6]
  assign _T_268 = _T_266 + _T_267; // @[VecMul.scala 42:21:@124.6]
  assign _T_269 = _T_266 + _T_267; // @[VecMul.scala 42:21:@125.6]
  assign _T_270 = io_A_11 * io_B_13; // @[VecMul.scala 42:35:@126.6]
  assign _T_271 = _T_269 + _T_270; // @[VecMul.scala 42:21:@127.6]
  assign ans_9 = _T_269 + _T_270; // @[VecMul.scala 42:21:@128.6]
  assign _T_273 = io_A_8 * io_B_2; // @[VecMul.scala 42:35:@129.6]
  assign _T_274 = {{1'd0}, _T_273}; // @[VecMul.scala 42:21:@130.6]
  assign _T_275 = _T_274[31:0]; // @[VecMul.scala 42:21:@131.6]
  assign _T_276 = io_A_9 * io_B_6; // @[VecMul.scala 42:35:@132.6]
  assign _T_277 = _T_275 + _T_276; // @[VecMul.scala 42:21:@133.6]
  assign _T_278 = _T_275 + _T_276; // @[VecMul.scala 42:21:@134.6]
  assign _T_279 = io_A_10 * io_B_10; // @[VecMul.scala 42:35:@135.6]
  assign _T_280 = _T_278 + _T_279; // @[VecMul.scala 42:21:@136.6]
  assign _T_281 = _T_278 + _T_279; // @[VecMul.scala 42:21:@137.6]
  assign _T_282 = io_A_11 * io_B_14; // @[VecMul.scala 42:35:@138.6]
  assign _T_283 = _T_281 + _T_282; // @[VecMul.scala 42:21:@139.6]
  assign ans_10 = _T_281 + _T_282; // @[VecMul.scala 42:21:@140.6]
  assign _T_285 = io_A_8 * io_B_3; // @[VecMul.scala 42:35:@141.6]
  assign _T_286 = {{1'd0}, _T_285}; // @[VecMul.scala 42:21:@142.6]
  assign _T_287 = _T_286[31:0]; // @[VecMul.scala 42:21:@143.6]
  assign _T_288 = io_A_9 * io_B_7; // @[VecMul.scala 42:35:@144.6]
  assign _T_289 = _T_287 + _T_288; // @[VecMul.scala 42:21:@145.6]
  assign _T_290 = _T_287 + _T_288; // @[VecMul.scala 42:21:@146.6]
  assign _T_291 = io_A_10 * io_B_11; // @[VecMul.scala 42:35:@147.6]
  assign _T_292 = _T_290 + _T_291; // @[VecMul.scala 42:21:@148.6]
  assign _T_293 = _T_290 + _T_291; // @[VecMul.scala 42:21:@149.6]
  assign _T_294 = io_A_11 * io_B_15; // @[VecMul.scala 42:35:@150.6]
  assign _T_295 = _T_293 + _T_294; // @[VecMul.scala 42:21:@151.6]
  assign ans_11 = _T_293 + _T_294; // @[VecMul.scala 42:21:@152.6]
  assign _T_297 = io_A_12 * io_B_0; // @[VecMul.scala 42:35:@153.6]
  assign _T_298 = {{1'd0}, _T_297}; // @[VecMul.scala 42:21:@154.6]
  assign _T_299 = _T_298[31:0]; // @[VecMul.scala 42:21:@155.6]
  assign _T_300 = io_A_13 * io_B_4; // @[VecMul.scala 42:35:@156.6]
  assign _T_301 = _T_299 + _T_300; // @[VecMul.scala 42:21:@157.6]
  assign _T_302 = _T_299 + _T_300; // @[VecMul.scala 42:21:@158.6]
  assign _T_303 = io_A_14 * io_B_8; // @[VecMul.scala 42:35:@159.6]
  assign _T_304 = _T_302 + _T_303; // @[VecMul.scala 42:21:@160.6]
  assign _T_305 = _T_302 + _T_303; // @[VecMul.scala 42:21:@161.6]
  assign _T_306 = io_A_15 * io_B_12; // @[VecMul.scala 42:35:@162.6]
  assign _T_307 = _T_305 + _T_306; // @[VecMul.scala 42:21:@163.6]
  assign ans_12 = _T_305 + _T_306; // @[VecMul.scala 42:21:@164.6]
  assign _T_309 = io_A_12 * io_B_1; // @[VecMul.scala 42:35:@165.6]
  assign _T_310 = {{1'd0}, _T_309}; // @[VecMul.scala 42:21:@166.6]
  assign _T_311 = _T_310[31:0]; // @[VecMul.scala 42:21:@167.6]
  assign _T_312 = io_A_13 * io_B_5; // @[VecMul.scala 42:35:@168.6]
  assign _T_313 = _T_311 + _T_312; // @[VecMul.scala 42:21:@169.6]
  assign _T_314 = _T_311 + _T_312; // @[VecMul.scala 42:21:@170.6]
  assign _T_315 = io_A_14 * io_B_9; // @[VecMul.scala 42:35:@171.6]
  assign _T_316 = _T_314 + _T_315; // @[VecMul.scala 42:21:@172.6]
  assign _T_317 = _T_314 + _T_315; // @[VecMul.scala 42:21:@173.6]
  assign _T_318 = io_A_15 * io_B_13; // @[VecMul.scala 42:35:@174.6]
  assign _T_319 = _T_317 + _T_318; // @[VecMul.scala 42:21:@175.6]
  assign ans_13 = _T_317 + _T_318; // @[VecMul.scala 42:21:@176.6]
  assign _T_321 = io_A_12 * io_B_2; // @[VecMul.scala 42:35:@177.6]
  assign _T_322 = {{1'd0}, _T_321}; // @[VecMul.scala 42:21:@178.6]
  assign _T_323 = _T_322[31:0]; // @[VecMul.scala 42:21:@179.6]
  assign _T_324 = io_A_13 * io_B_6; // @[VecMul.scala 42:35:@180.6]
  assign _T_325 = _T_323 + _T_324; // @[VecMul.scala 42:21:@181.6]
  assign _T_326 = _T_323 + _T_324; // @[VecMul.scala 42:21:@182.6]
  assign _T_327 = io_A_14 * io_B_10; // @[VecMul.scala 42:35:@183.6]
  assign _T_328 = _T_326 + _T_327; // @[VecMul.scala 42:21:@184.6]
  assign _T_329 = _T_326 + _T_327; // @[VecMul.scala 42:21:@185.6]
  assign _T_330 = io_A_15 * io_B_14; // @[VecMul.scala 42:35:@186.6]
  assign _T_331 = _T_329 + _T_330; // @[VecMul.scala 42:21:@187.6]
  assign ans_14 = _T_329 + _T_330; // @[VecMul.scala 42:21:@188.6]
  assign _T_333 = io_A_12 * io_B_3; // @[VecMul.scala 42:35:@189.6]
  assign _T_334 = {{1'd0}, _T_333}; // @[VecMul.scala 42:21:@190.6]
  assign _T_335 = _T_334[31:0]; // @[VecMul.scala 42:21:@191.6]
  assign _T_336 = io_A_13 * io_B_7; // @[VecMul.scala 42:35:@192.6]
  assign _T_337 = _T_335 + _T_336; // @[VecMul.scala 42:21:@193.6]
  assign _T_338 = _T_335 + _T_336; // @[VecMul.scala 42:21:@194.6]
  assign _T_339 = io_A_14 * io_B_11; // @[VecMul.scala 42:35:@195.6]
  assign _T_340 = _T_338 + _T_339; // @[VecMul.scala 42:21:@196.6]
  assign _T_341 = _T_338 + _T_339; // @[VecMul.scala 42:21:@197.6]
  assign _T_342 = io_A_15 * io_B_15; // @[VecMul.scala 42:35:@198.6]
  assign _T_343 = _T_341 + _T_342; // @[VecMul.scala 42:21:@199.6]
  assign ans_15 = _T_341 + _T_342; // @[VecMul.scala 42:21:@200.6]
  assign io_C_0 = ans_0[15:0]; // @[VecMul.scala 51:8:@223.4]
  assign io_C_1 = ans_1[15:0]; // @[VecMul.scala 51:8:@224.4]
  assign io_C_2 = ans_2[15:0]; // @[VecMul.scala 51:8:@225.4]
  assign io_C_3 = ans_3[15:0]; // @[VecMul.scala 51:8:@226.4]
  assign io_C_4 = ans_4[15:0]; // @[VecMul.scala 51:8:@227.4]
  assign io_C_5 = ans_5[15:0]; // @[VecMul.scala 51:8:@228.4]
  assign io_C_6 = ans_6[15:0]; // @[VecMul.scala 51:8:@229.4]
  assign io_C_7 = ans_7[15:0]; // @[VecMul.scala 51:8:@230.4]
  assign io_C_8 = ans_8[15:0]; // @[VecMul.scala 51:8:@231.4]
  assign io_C_9 = ans_9[15:0]; // @[VecMul.scala 51:8:@232.4]
  assign io_C_10 = ans_10[15:0]; // @[VecMul.scala 51:8:@233.4]
  assign io_C_11 = ans_11[15:0]; // @[VecMul.scala 51:8:@234.4]
  assign io_C_12 = ans_12[15:0]; // @[VecMul.scala 51:8:@235.4]
  assign io_C_13 = ans_13[15:0]; // @[VecMul.scala 51:8:@236.4]
  assign io_C_14 = ans_14[15:0]; // @[VecMul.scala 51:8:@237.4]
  assign io_C_15 = ans_15[15:0]; // @[VecMul.scala 51:8:@238.4]
  assign io_valid = io_load; // @[VecMul.scala 47:14:@201.6 VecMul.scala 49:14:@204.6]
endmodule
